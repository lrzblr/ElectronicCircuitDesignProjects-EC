* deney 7


VGS 4 0 0V
VDS 6 0 0V

R1 3 6 1k



M1 3 2 0 0 N3306M
RG 4 2 270
RL 3 0 1.2E8
C1 2 0 28E-12
C2 3 2 3E-12 
D1 0 3 N3306D
.MODEL N3306M NMOS VTO=1.824 RS=1.572 RD=1.436 IS=1E-15 KP=.1233
+CBD=35E-12 PB=1
.MODEL N3306D D IS=5E-12 RS=.768


 .DC VDS 0 10 0.5 VGS  0 2 0.5 
 .PROBE
 .END