*C51
Vi 4 0 sin(0 20mV 1khz)
VCC 1 0 DC 12V
Q1 5 2 10 BC547B
Q2 7 6 9 BC547B
C1b 2 3 10uF
C1e 10 11 100uF
C2 5 6 10uF
C2e 9 0 100uF
C22 7 8 10uF
c23 8 12 10uF
R21 3 4 180k
R22 3 0 20k
R23 2 0 22k
R11 1 2 68k
R1c 1 5 4.7k
R6 10 11 2.2k
R52 11 0 100
R111 1 6 47k
R24 6 0 33k
R51 1 7 2.2k
R11e 9 0 2.2k
R12l 8 0 1k
R2f 11 12 4.7k
.MODEL BC547B NPN BF=500 NE=1.3 ISE=9.72F IKF=80M IS=20F VAF=50 +ikr=12m BR=10 NC=2 VAR=10 RB=280 RE=1 RC=40 VJE=.48 tr=.3u tf=.5n +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc=.33 isc=47p kf=2f
.PROBE
.TRAN 1us 4ms
.END