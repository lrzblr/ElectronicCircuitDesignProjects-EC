*C63
VCC 1 0 DC 12V
Vi 3 0 sin(0 20mV 1khz)
Q1 4 2 6 BC547B
R1 1 2 68k
R2 2 0 15k
R4 1 4 4.7k
R5 6 0 1.2k
Rload 5 0 1k
Cb1 2 3 22uF
Cb2 4 5 22uF
Ce 6 0 47uF
*sekil7 icin
rf 2 7 47k
cf 7 4 22uF
.MODEL BC547B NPN BF=500 NE=1.3 ISE=9.72F IKF=80M IS=20F VAF=50 +ikr=12m BR=10 NC=2 VAR=10 RB=280 RE=1 RC=40 VJE=.48 tr=.3u tf=.5n +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc=.33 isc=47p kf=2f
.PROBE
.TRAN 1us 5ms
.END