*
VDC 1 0 DC 12V
Vi 3 0 sin(0 200mV 1khz)
R1 1 2 110k
R2 2 0 10k
R3 1 4 1.5k
R4 7 0 24
R5 1 8 120
R6 10 0 120
Rload 11 0 1.2k
C1 2 3 1uF
C2 9 11 1uF
Q1 6 2 7 BD135
Q2 8 4 9 BD135
Q3 9 6 10 BD136
D1 4 5 1N4001
D2 5 6 1N4001
.model 1N4001 D(Is=14.11n N=1.984 Rs=33.89m Ikf=94.81 Xti=3 Eg=1.11 Cjo=25.89p M=.44 Vj=.3245 Fc=.5 Bv=75 Ibv=10u Tt=5.7u Iave=1 Vpk=50 mfg=GI type=silicon)
.model BD135 NPN(Is=40f Xti=3 Eg=1.11 Vaf=115.7 Bf=180.2 Ise=40f Ne=1.363 Ikf=4.927 Nk=1.247 Xtb=1.5 Br=10 Isc=85f Nc=2 Ikr=0 Rc=0 Cjc=19.23p Mjc=.3439 Vjc=.5635 Fc=.5 Cje=60.49p Mje=.3589 Vje=.7585 Tr=116n Tf=550p Itf=1 Xtf=0 Vtf=10 QCO=1E-10 GAMMA=1E-8 RCO=5)
.model BD136 PNP (Is=10f Xti=3 Eg=1.11 Vaf=95.7 Bf=178.7 Ise=134.1f Ne=1.553 Ikf=2 Nk=.8366 Xtb=1.5 Br=5 Isc=85f Nc=2 Ikr=0 Rc=0 Cjc=60p Mjc=.4 Vjc=.8 Fc=.8 Cje=115.6p Mje=.3766 Vje=.7703 Tr=116n Tf=500p Itf=1 Xtf=0 Vtf=10 QCO=1E-10 GAMMA=5n RCO=5)
.PROBE
.TRAN 1us 5ms
.END