*deney3

R1 2 3 120k
R2 1 4 1k
Vcc 1 0 DC 0.2V 
Vbb 2 0 DC 1V 
Q1 4 3  0 BC237
.MODEL BC237 NPN IS =1.8E-14 ISE=5.0E-14 NF =.9955 NE =1.46 BF =400 BR =35.5 IKF=.14 IKR=.03 ISC=1.72E-13 NC =1.27 NR =1.005 RB =.56 RE =.6 RC =.25 VAF=80 VAR=12.5 CJE=13E12 TF =.64E-9 CJC=4E-12 TR =50.72E-9 VJC=.54 MJC=.33 
.DC Vcc LIST 0.2, 1, 3, 5, 7, 9, 11, 13, 15 Vbb LIST 0.1 0.2 0.3 0.4 0.5 0.6 0.7  0.8 0.9 1
.probe
.end