*

VCC 1 0 12V
VEE 0 3 12V
V1 5 0 sin(0 10mV 1kHz)
V2 8 0 0
R1 1 2 10K
R3 1 4 10K
R4 1 7 10K
M1 4 5 6 3 BS170
M2 7 8 6 3 BS170
M3 6 2 3 3 BS170
M4 2 2 3 3 BS170
.MODEL BS170 NMOS VTO=1.824 RS=1.572 RD=1.436 IS=1E-15 KP=.1233 CBD=35E-12 PB=1
.PROBE
.TRAN 1US