*C71
Vi 7 0 sin(0 1V 1khz)
Vcc_p 1 0 DC 12V
Vcc_n 6 0 DC -12V
R1 1 2 120
R2 5 6 120
R3 8 0 1.2k
C1 3 7 1uF
C2 4 8 1uF
Q1 2 3 4 BC547B
Q2 4 3 5 BD136
.MODEL BC237 NPN IS =1.8E-14 ISE=5.0E-14 NF =.9955 NE =1.46 BF =400 BR =35.5 IKF=.14 IKR=.03 ISC=1.72E-13 NC =1.27 NR =1.005 RB =.56 RE =.6 RC =.25 VAF=80 VAR=12.5 CJE=13E-12 TF =.64E-9 CJC=4E-12 TR =50.72E-9 VJC=.54 MJC=.33
Teslim Tarihi: 26 Nisan 2022 10.00
**.MODEL BD135 NPN IC_VBE=1.10250E-36 IC_VCE=1.10250E-36 STATE=1 TEMP=0 AREA=1.0 STATE_FACTOR=0 IS=90.36e-9 BF=95. NF=2.03 VAF=200 IKF=500.0 ISE=1.039e-6 NE=17.89 BR=8.423 NR=2.03 VAR=10.0 ISC=0 NC=1 RB=0.9454 RBM=0.9454 RE=0.01 RC=0.3758 CJE=100.0e-12 VJE=0.7 MJE=0.4 TF=568.41e-12 XTF=0 ITF=0 CJC=100e-12 VJC=0.7 MJC=0.4 XCJC=0.500 CJS=0 XTB=1.5
**.MODEL BD136 PNP IC_VCE=1.10250E-36 IC_VBE=1.10250E-36 STATE=1 TEMP=0 AREA=1 STATE_FACTOR=0 IS=2.900E-13 BF=1.237E+02 NF=1.079E+00 VAF=1.000E+02 IKF=4.474E-01 ISE=7.453E-12 NE=1.820E+00 BR=3.434E-01 NR=1.181E+00 VAR=5.000E+01 IKR=1.000E+09 ISC=0.000E+00 NC=2.000E+00 RB=3.700E-01 IRB=1.500E-01 RBM=3.700E-01 RE=9.600E-02 RC=5.520E-01 CJE=2.100E-10 VJE=7.500E-01 MJE=3.300E-01 TF=1.853E-09 XTF=8.483E-01 VTF=9.990E+05 ITF=1.696E+00 PTF=0.000E+00 CJC=1.000E-10 VJC=7.500E-01 MJC=3.300E-01 XCJC=1.000E+00 TR=0.000E+00 CJS=1.000E-12 VJS=7.500E-01 MJS=0.000E+00 XTB=1.500E+00 EG=1.110E+00 XTI=1.000E+00 FC=5.000E-01
.MODEL BD136 PNP(Is=10f Xti=3 Eg=1.11 Vaf=95.7 Bf=178.7 Ise=134.1f Ne=1.553 Ikf=2 Nk=.8366 Xtb=1.5 Br=5 Isc=85f Nc=2 Ikr=0 Rc=0 Cjc=60p Mjc=.4 Vjc=.8 Fc=.8 Cje=115.6p Mje=.3766 Vje=.7703 Tr=116n Tf=500p Itf=1 Xtf=0 Vtf=10 QCO=1E-10 GAMMA=5n RCO=5)
.PROBE
.TRAN 1us 5ms
.END