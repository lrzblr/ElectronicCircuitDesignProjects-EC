*
VCC 1 0 DC 12V
Vi 3 0 sin(0 110mV 1khz)
R1 1 2 110k
R2 1 4 1.5k
R3 2 0 10k
R4 5 0 24
R5 6 0 2.2k
C1 2 3 1uF
C2 4 6 1uF
Q1 4 2 5 BC237
.MODEL BC237 NPN IS =1.8E-14 ISE=5.0E-14 NF =.9955 NE =1.46 BF =400 BR =35.5 IKF=.14 IKR=.03 ISC=1.72E-13 NC =1.27 NR =1.005 RB =.56 RE =.6 RC =.25 VAF=80 VAR=12.5 CJE=13E-12 TF =.64E-9 CJC=4E-12 TR =50.72E-9 VJC=.54 MJC=.33
.PROBE
.TRAN 1us 5ms
.END