*deney9.1


VCC 5 0 12V
Vs 1 0 sin(0 20mV 1kHz)

C1 2 1 1u
C2 4 6 1u
C3 7 9 1u

RB2 2 0 10k
RB1 2 5 100k
RC1 5 4 2.2k
RE1 3 0 270
RB3 5 6 100k
RB4 6 0 10k
RC2 5 7 2.2k
RE2 8 0 1k
R5 9 0 1T

Q1 4 2 3 BC237
Q2 7 6 8 BC237

.MODEL BC237 NPN IS =1.8E-14 ISE=5.0E-14 NF =.9955 NE =1.46 BF =400 BR =35.5 IKF=.14 IKR=.03 ISC=1.72E-13 NC =1.27 NR =1.005 RB =.56 RE =.6 RC =.25 VAF=80 VAR=12.5 CJE=13E-12 TF =.64E-9 CJC=4E-12 TR =50.72E-9 VJC=.54 MJC=.33

.PROBE 
.TRAN 0ms 2ms 0.001ms
.END
