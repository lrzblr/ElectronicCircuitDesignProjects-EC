**
V1 1 0 AC 20mV
V2 3 0 DC 12V
Cs 2 1 10uF
R1 3 2 82K
R2 2 0 8.2K
Rc 3 4 12K
Cc 4 0 470uF
Q1 4 2 5 BC237
RE 5 0 1K
Ce 5 6 10uF
Rl 6 0 3.3K
C4 6 0 1nF
.MODEL BC237 NPN IS =1.8E-14 ISE=5.0E-14 NF =.9955 NE =1.46 BF =400 BR =35.5 IKF=.14 IKR=.03 ISC=1.72E-13 NC =1.27 NR=1.005 RB =.56 RE =.6 RC =.25
VAF=80 VAR=12.5 CJE=13E-12 TF =.64E-9 CJC=4E-12 TR =50.72E-9 VJC=.54 MJC=.33
.AC DEC 10 1HZ 100MEG
.PROBE
.END