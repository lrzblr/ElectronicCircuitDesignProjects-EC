* deney4

Vg 1 0 PULSE(0 9 2 0 0 2 4)
R1 1 2 100k
R2  2 3 100k
R3 3 6 1k
R4 4 5 330
C1 3 0 220u
D1 1 4 LED
Q1 5  6  0 BC237



.model LED D (IS=93.2P RS=42M N=3.73 BV=4 IBV=10U  CJO=2.97P VJ=.75 M=.333 TT=4.32U)
.MODEL BC237 NPN IS =1.8E-14 ISE=5.0E-14 NF =.9955 NE =1.46 BF =400 BR =35.5 IKF=.14 IKR=.03 ISC=1.72E-13 NC =1.27 NR =1.005 RB =.56 RE =.6 RC =.25 VAF=80 VAR=12.5 CJE=13E-12 TF =.64E-9 CJC=4E-12 TR =50.72E-9 VJC=.54 MJC=.33
.TRAN 1ms 16s 
.PROBE
.END