*
.param Rval 10k
V1 1 0 12V
R1 1 2 1K
R2 1 4 1K
R3 2 3 {Rval}
.STEP PARAM Rval 1K 10K 1K
M1 3 3 0 BS170
M2 4 3 0 BS170
.MODEL BS170 NMOS VTO=1.824 RS=1.572 RD=1.436 IS=1E-15 KP=.1233 CBD=35E-12 PB=1
.OP .TRAN 0 100ns 0
.PROBE
.END