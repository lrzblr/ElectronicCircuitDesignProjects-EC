**
V1 6 0 AC 20mV;
V2 3 0 DC 12V;
R1 4 0 360k;
R2 1 0 220;
R3 3 4 1M;
R4 3 2 1k;
R5 5 0 10k;
C1 4 6 1uF;
C2 1 0 1uF;
C3 2 5 1uF;
M1 3 2 0 0 N3306M
RG 4 2 270
RL 3 0 1.2E8
C1 2 0 28E-12
C2 3 2 3E-12
D1 0 3 N3306D
.MODEL N3306M NMOS VTO=1.824 RS=1.572 RD=1.436 IS=1E-15 KP=.1233
+CBD=35E-12 PB=1
.MODEL N3306D D IS=5E-12 RS=.768
.AC dec 10 1Hz 100000kHz;
.probe;