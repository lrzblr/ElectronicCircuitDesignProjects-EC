*
.param Rval 10k
V1 1 0 12V
R1 1 2 1k
R2 1 4 1k
R3 2 3 {Rval}
.step param Rval 1k 10k 1k
Q1 3 3 0 BC237
Q2 4 3 0 BC237
.model BC237 NPN IS =1.8E-14 ISE=5.0E-14 NF =.9955 NE =1.46 BF =400 BR =35.5 IKF=.14 IKR=.03 ISC=1.72E-13 NC =1.27 NR =1.005 RB =.56 RE =.6 RC =.25 VAF=80 VAR=12.5 CJE=13E-12 TF =.64E-9 CJC=4E-12 TR =50.72E-9 VJC=.54 MJC=.33
.op
.tran 0 100ns 0
.probe
.end