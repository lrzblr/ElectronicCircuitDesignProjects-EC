*deney 2

V1 1 0 sin(0 6V 50hz)
V2 2 1 sin(0 6V 50hz)

C1 5 3 100U
R1 5 3 100K

D1 3 2 D1N4001
D2 3 0 D1N4001
D3 2 5 D1N4001
D4 0 5 D1N4001

.MODEL D1N4001 D(Is=14.11n N=1.984 Rs=33.89m Ikf=94.81 Xti=3 Eg=1.11 Cjo=25.89p M=.44 Vj=.3245 Fc=.5 Bv=75 Ibv=10u Tt=5.7u)
.PROBE 
.TRAN 0.1ms 40ms 0.1ms
 .END

