*
Vi1 1 0 sin(0 10m 1khz)
Vi2 7 0 DC 0V
V3 4 0 DC 12V
V4 0 9 DC 12V
R1 1 2 1k
R2 7 6 1k
R3 3 4 10k
R4 4 5 10k
R5 4 10 22k
Q1 3 2 8 BC237
Q2 5 6 8 BC237
Q3 8 10 9 BC237
Q4 10 10 9 BC237
.MODEL BC237 NPN IS =1.8E-14 ISE=5.0E-14 NF =.9955 NE =1.46 BF =400 BR =35.5 IKF=.14 IKR=.03 ISC=1.72E-13 NC =1.27 NR =1.005 RB =.56 RE =.6 RC =.25 VAF=80 VAR=12.5 CJE=13E-12 TF =.64E-9 CJC=4E-12 TR =50.72E-9 VJC=.54 MJC=.33
.TRAN 0.1ms 4ms
.PROBE
.END